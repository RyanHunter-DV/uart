
// register address & name
parameter DRAddr = 10'h0;

// RSR receive status register, RO
parameter RSRAddr = 10'h1;
// ECR Error clear, WO
parameter ECRAddr=10'h1;
... //TODO, require more